LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;
USE ieee.Numeric_Std.ALL;

ENTITY mikroMemory IS
	PORT (
		addr : IN STD_LOGIC_VECTOR(7 DOWNTO 0); -- address
		dat_out  : OUT STD_LOGIC_VECTOR(76 DOWNTO 0); -- data to write
		clk : IN STD_LOGIC -- clock
	);
END ENTITY mikroMemory;

ARCHITECTURE description OF mikroMemory IS

   TYPE ram_type IS ARRAY (0 TO 159) OF STD_LOGIC_VECTOR(76 DOWNTO 0);
   SIGNAL ram : ram_type;

BEGIN	
	dat_out <= ram(to_integer(unsigned(addr)));


	ram(0) <= "00001110000000000000000000000000000000000000000000000000000000000000000000000";
	ram(1) <= "00000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(2) <= "00000000000000000000000000000000000000000000000000000000010000001100000000000";
	ram(3) <= "10000000001000000000000000000000000000000000000000000000000000000000000000000";
	ram(4) <= "00000000000000000000000000000000000000000000000000000000000000000000000000100";
	ram(5) <= "01000000000010000000000000000000000000000000000000000000000000000000000000000";
	ram(6) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(7) <= "00000001000000000000000000000000000000000000000000000000000000000000000000000";
	ram(8) <= "00000000000000000000000000000000000000000000000000000000000000000000100001111";
	ram(9) <= "01000000000010000000000000000000000000000000000000000000000000000000000000000";
	ram(10) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(11) <= "00000000100000000000000000000000000000000000000000000000000000000001000001111";
	ram(12) <= "01000000000010000000000000000000000000000000000000000000000000000000000000000";
	ram(13) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(14) <= "00000000010000000000000000000000000000000000000000000000000000000000000000000";
	ram(15) <= "00000000000000000000000000000000000000000000000000000000000000001011100000000";
	ram(16) <= "00000000000001000000000000000000000000000000000000000000000000000001110001001";
	ram(17) <= "00000000000000000000000000000000000000000000000000000000000000000001110001001";
	ram(18) <= "01100000000000000001000000000000000000000000000000000000000000000000000000000";
	ram(19) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(20) <= "01100000000000100001000000000000000000000000000000000000000000000000000000000";
	ram(21) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(22) <= "00000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(23) <= "00000000000000000000010000000000000000000000000000000000000000000000000000000";
	ram(24) <= "01100000000000000001000000000000000000000000000000000000000000000000000000000";
	ram(25) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(26) <= "01100000000000100001000000000000000000000000000000000000000000000000000000000";
	ram(27) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(28) <= "00000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(29) <= "00000000001000000000000000000000000000000000000000000000000000000001110001001";
	ram(30) <= "00000000000000000000001000000000000000000000000000000000000000000001110001001";
	ram(31) <= "00000000000000000000000100000000000000000000000000000000000000000001110001001";
	ram(32) <= "00000000000000000000000010000000000000000000000000000000000000000001110001001";
	ram(33) <= "00000000000000000000000001000000000000000000000000000000000000000001110001001";
	ram(34) <= "00000000000000000000000000000000000000000000000000000000000000000010010001001";
	ram(35) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(36) <= "00000000000000000000000000000000000000000000000000000000000000000010110001001";
	ram(37) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(38) <= "00000000000000000000000000000000000000000000000000000000000000000011010001001";
	ram(39) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(40) <= "00000000000000000000000000000000000000000000000000000000000000000011110001001";
	ram(41) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(42) <= "00000000000000000000000000000000000000000000000000000000000000000100010001001";
	ram(43) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(44) <= "00000000000000000000000000000000000000000000000000000000000000000100110001001";
	ram(45) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(46) <= "00000000000000000000000000000000000000000000000000000000000000000101010001001";
	ram(47) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(48) <= "00000000000000000000000000000000000000000000000000000000000000000101110001001";
	ram(49) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(50) <= "00000000000000000000000000000000000000000000000000000000000000000110010001001";
	ram(51) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(52) <= "00000000000000000000000000000000000000000000000000000000000000000110110001001";
	ram(53) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(54) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(55) <= "00000000000000000000000000000100000000000000000000000000000000000000000000000";
	ram(56) <= "00000000000000000000000000000000000000000000000000000000000000000111010001001";
	ram(57) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(58) <= "00000000000000000000000000000100000000000000000000000000000000000000000000000";
	ram(59) <= "00000000000000000000000000000000000000000000000000000000000000000111110001001";
	ram(60) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(61) <= "00000000000000000000000000000100000000000000000000000000000000000000000000000";
	ram(62) <= "00000000000000000000000000000000000000000000000000000000000000001000010001001";
	ram(63) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(64) <= "00000000000000110010100000000000000000000000000000000000000000000000000000000";
	ram(65) <= "01101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(66) <= "00000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(67) <= "01101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(68) <= "00000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(69) <= "00000000001100000000000000101000000000000000000000000000000000000001110001001";
	ram(70) <= "00000000000000110010100000000000000000000000000000000000000000000000000000000";
	ram(71) <= "01101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(72) <= "00000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(73) <= "01101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(74) <= "00000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(75) <= "00000000000000110100100000000000000000000000000000000000000000000000000000000";
	ram(76) <= "01101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(77) <= "00000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(78) <= "01101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(79) <= "00000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(80) <= "00000000001100000000001000101000000000000000000000000000000000000001100000100";
	ram(81) <= "00000000000000000000000000000000111000111000000000000000000000000001110001001";
	ram(82) <= "00000000000000000000000000000000101000111000000000000000000000000001110001001";
	ram(83) <= "00000000000000000000000000000000000001111000000000000000000000000001110001001";
	ram(84) <= "00000000000000000000000000000000001001111000000000000000000000000001110001001";
	ram(85) <= "00000000000000000000000000000001001010111000000000000000000000000001110001001";
	ram(86) <= "00000000000000000000000000000001010010111000000000000000000000000001110001001";
	ram(87) <= "00000000000000000000000000000001001100111000000000000000000000000001110001001";
	ram(88) <= "00000000000000000000000000000001010011111000000000000000000000000001110001001";
	ram(89) <= "00000000000000000000000000000000000000000000000000000000000000000001110001001";
	ram(90) <= "00000000000000000000000000000001010100111000000000000000000000000001110001001";
	ram(91) <= "00000000000000000000000000000001001000111000000000000000000000000001110001001";
	ram(92) <= "00000000000000000000000000000001010000111000000000000000000000000001110001001";
	ram(93) <= "01100000000000000001000000000000000000000000000000000000000000000000000000000";
	ram(94) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(95) <= "01100000000000100001000000000000000000000000000000000000000000000000000000000";
	ram(96) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(97) <= "00000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(98) <= "00000000000000000000000000000000000000100000000000000000000000000001110001001";
	ram(99) <= "00000000000000110000100000000000000000000000000001000000000000000000000000000";
	ram(100) <= "01101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(101) <= "00000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(102) <= "01101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(103) <= "00000000000000000000000000000010000000000000000000000000000000000001110001001";
	ram(104) <= "00000000000000000000000000000000000000111000000000000000000000000001110001001";
	ram(105) <= "00000000000000000000000000000000001000111000000000000000000000000001110001001";
	ram(106) <= "00000000000000000000000000000001011000111000000000000000000000000001110001001";
	ram(107) <= "00000000000000000000000000000000010000111000000000000000000000000001110001001";
	ram(108) <= "00000000000000000000000000000000011000111000000000000000000000000001110001001";
	ram(109) <= "00000000000000000000000000000000100000111000000000000000000000000001110001001";
	ram(110) <= "00000000000000000000000000000000001000010000000000000000000000000001110001001";
	ram(111) <= "00000000000000000000000000000000010000010000000000000000000000000001110001001";
	ram(112) <= "00000000000000000000000000000000000000000000000000000000000000001000110001000";
	ram(113) <= "00000000000000000000000000000000000000000111000000000000000000000000000000000";
	ram(114) <= "00000000000000000000000000000000001000010000011010000000000000000000000000000";
	ram(115) <= "00000000000000000000000000000000000000000000000000000000000000001001001110010";
	ram(116) <= "00000000000000000000000000000000000000000000101010000000000000000000000000000";
	ram(117) <= "00000000000000000000000000000000000000000110001110000000000000000001110001001";
	ram(118) <= "00000000000000111110000000000000000000000000000000000000000000000000000000000";
	ram(119) <= "00000000000000000000000000000000000000100000000000000000000000000001110001001";
	ram(120) <= "01010000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(121) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(122) <= "00000000000000100000000000000000000000000000000000000000010000000000000000000";
	ram(123) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(124) <= "00000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(125) <= "00000000000000000000000000000000000000100000000000000000000000000001110001001";
	ram(126) <= "01010000000000110000000000000000000000000000000001000000000000000000000000000";
	ram(127) <= "00001010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(128) <= "00000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(129) <= "00001100000000000000000000000000000000000000000000000000010000000000000000000";
	ram(130) <= "00000000000000000000000000000010000000000000000000000000000000000001110001001";
	ram(131) <= "00000000000000000000000000000000110000101000000000000000000000000000000000000";
	ram(132) <= "00000000000000000000000000000000101000101000000000000000000000000001110001001";
	ram(133) <= "00000000000000000000000000000000000000000000001100000000000000000001110001001";
	ram(134) <= "00000000000000000000000000000000000000000000000000100000000000000001110001001";
	ram(135) <= "00000000000000000000000000000000000000000000000000010000000000000001110001001";
	ram(136) <= "00000000000000000000000000000000000000000000000000001000000000000000000000000";
	ram(137) <= "00000000000000000000000000000000000000000000000000000000000000001001110001011";
	ram(138) <= "00000000000000000000000000000000000000000000000000000110101000000001110010001";
	ram(139) <= "00000000000000000000000000000000000000000000000000000000000000001010010001101";
	ram(140) <= "00000000000000000000000000000000000000000000000000000111000100000001110010001";
	ram(141) <= "00000000000000000000000000000000000000000000000000000000000000001010110001111";
	ram(142) <= "00000000000000000000000000000000000000000000000000000111100010000001110010001";
	ram(143) <= "00000000000000000000000000000000000000000000000000000000000000001011000000100";
	ram(144) <= "00000000000000000000000000000000000000000000000000000100000000000000000000000";
	ram(145) <= "00000000000000110010100000000000000000000000000000000000000000000000000000000";
	ram(146) <= "01101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(147) <= "00000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(148) <= "01101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(149) <= "00000000000000110100100000000010000000000000000000000000000000000000000000000";
	ram(150) <= "01101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(151) <= "00000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(152) <= "01101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(153) <= "00000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(154) <= "01110000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(155) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(156) <= "00000000000000100000000000000000000000000000000000000000010000000000000000000";
	ram(157) <= "00001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(158) <= "00000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(159) <= "00000000001000000000001000000000000000000000000000000000000000000001100000100";



	
END description;



--00 00 00 00 00 00 00 00		00 00
