LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;
USE ieee.Numeric_Std.ALL;

ENTITY mikroMemory IS
	PORT (
		addr : IN STD_LOGIC_VECTOR(7 DOWNTO 0); -- address
		dat_out  : OUT STD_LOGIC_VECTOR(75 DOWNTO 0); -- data to write
		clk : IN STD_LOGIC -- clock
	);
END ENTITY mikroMemory;

ARCHITECTURE description OF mikroMemory IS

   TYPE ram_type IS ARRAY (0 TO 157) OF STD_LOGIC_VECTOR(75 DOWNTO 0);
   SIGNAL ram : ram_type;

BEGIN	
	dat_out <= ram(to_integer(unsigned(addr)));

	ram(0) <= "0000000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(1) <= "1000000000010000000000000000000000000000000000000000000000000000000000000000";
	ram(2) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(3) <= "0000001000000000000000000000000000000000000000000000000000000000000000000000";
	ram(4) <= "0000000000000000000000000000000000000000000000000000000000000000000100001011";
	ram(5) <= "1000000000010000000000000000000000000000000000000000000000000000000000000000";
	ram(6) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(7) <= "0000000100000000000000000000000000000000000000000000000000000000001000001011";
	ram(8) <= "1000000000010000000000000000000000000000000000000000000000000000000000000000";
	ram(9) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(10) <= "0000000010000000000000000000000000000000000000000000000000000000000000000000";
	ram(11) <= "0000000000000000000000000000000000000000000000000000000000000001011100000000";
	ram(12) <= "0000000000001000000000000000000000000000000000000000000000000000001110000101";
	ram(13) <= "0000000000000000000000000000000000000000000000000000000000000000001110000101";
	ram(14) <= "1100000000000000001000000000000000000000000000000000000000000000000000000000";
	ram(15) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(16) <= "1100000000000100001000000000000000000000000000000000000000000000000000000000";
	ram(17) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(18) <= "0000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(19) <= "0000000000000000000010000000000000000000000000000000000000000000000000000000";
	ram(20) <= "1100000000000000001000000000000000000000000000000000000000000000000000000000";
	ram(21) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(22) <= "1100000000000100001000000000000000000000000000000000000000000000000000000000";
	ram(23) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(24) <= "0000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(25) <= "0000000001000000000000000000000000000000000000000000000000000000001110000101";
	ram(26) <= "0000000000000000000001000000000000000000000000000000000000000000001110000101";
	ram(27) <= "0000000000000000000000100000000000000000000000000000000000000000001110000101";
	ram(28) <= "0000000000000000000000010000000000000000000000000000000000000000001110000101";
	ram(29) <= "0000000000000000000000001000000000000000000000000000000000000000001110000101";
	ram(30) <= "0000000000000000000000000000000000000000000000000000000000000000010110000101";
	ram(31) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(32) <= "0000000000000000000000000000000000000000000000000000000000000000010110000101";
	ram(33) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(34) <= "0000000000000000000000000000000000000000000000000000000000000000011110000101";
	ram(35) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(36) <= "0000000000000000000000000000000000000000000000000000000000000000011110000101";
	ram(37) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(38) <= "0000000000000000000000000000000000000000000000000000000000000000100010000101";
	ram(39) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(40) <= "0000000000000000000000000000000000000000000000000000000000000000100110000101";
	ram(41) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(42) <= "0000000000000000000000000000000000000000000000000000000000000000101110000101";
	ram(43) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(44) <= "0000000000000000000000000000000000000000000000000000000000000000101110000101";
	ram(45) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(46) <= "0000000000000000000000000000000000000000000000000000000000000000110110000101";
	ram(47) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(48) <= "0000000000000000000000000000000000000000000000000000000000000000110110000101";
	ram(49) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(50) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(51) <= "0000000000000000000000000000100000000000000000000000000000000000000000000000";
	ram(52) <= "0000000000000000000000000000000000000000000000000000000000000000111010000101";
	ram(53) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(54) <= "0000000000000000000000000000100000000000000000000000000000000000000000000000";
	ram(55) <= "0000000000000000000000000000000000000000000000000000000000000000111110000101";
	ram(56) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(57) <= "0000000000000000000000000000100000000000000000000000000000000000000000000000";
	ram(58) <= "0000000000000000000000000000000000000000000000000000000000000001000010000101";
	ram(59) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(60) <= "0000000000000110010100000000000000000000000000000000000000000000000000000000";
	ram(61) <= "1101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(62) <= "0000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(63) <= "1101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(64) <= "0000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(65) <= "0000000001100000000000000101000000000000000000000000000000000000001110000101";
	ram(66) <= "0000000000000110010100000000000000000000000000000000000000000000000000000000";
	ram(67) <= "1101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(68) <= "0000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(69) <= "1101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(70) <= "0000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(71) <= "0000000000000110100100000000000000000000000000000000000000000000000000000000";
	ram(72) <= "1101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(73) <= "0000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(74) <= "1101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(75) <= "0000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(76) <= "0000000001100000000000000101000000000000000000000000000000000000001100000000";
	ram(77) <= "0000000000000000000000000000000111000111000000000000000000000000001110000101";
	ram(78) <= "0000000000000000000000000000000101000111000000000000000000000000001110000101";
	ram(79) <= "0000000000000000000000000000000000001111000000000000000000000000001110000101";
	ram(80) <= "0000000000000000000000000000000001001111000000000000000000000000001110000101";
	ram(81) <= "0000000000000000000000000000001001010111000000000000000000000000001110000101";
	ram(82) <= "0000000000000000000000000000001010010111000000000000000000000000001110000101";
	ram(83) <= "0000000000000000000000000000001001100111000000000000000000000000001110000101";
	ram(84) <= "0000000000000000000000000000001010011111000000000000000000000000001110000101";
	ram(85) <= "0000000000000000000000000000000000000000000000000000000000000000001110000101";
	ram(86) <= "0000000000000000000000000000001010100111000000000000000000000000001110000101";
	ram(87) <= "0000000000000000000000000000001001000111000000000000000000000000001110000101";
	ram(88) <= "0000000000000000000000000000001010000111000000000000000000000000001110000101";
	ram(89) <= "1100000000000000001000000000000000000000000000000000000000000000000000000000";
	ram(90) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(91) <= "1100000000000100001000000000000000000000000000000000000000000000000000000000";
	ram(92) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(93) <= "0000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(94) <= "0000000000000000000000000000000000000100000000000000000000000000001110000101";
	ram(95) <= "0000000000000110000100000000000000000000000000001000000000000000000000000000";
	ram(96) <= "1101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(97) <= "0000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(98) <= "1101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(99) <= "0000000000000000000000000000010000000000000000000000000000000000001110000101";
	ram(100) <= "0000000000000000000000000000000000000110000000000000000000000000001110000101";
	ram(101) <= "0000000000000000000000000000000001000110000000000000000000000000001110000101";
	ram(102) <= "0000000000000000000000000000001011000110000000000000000000000000001110000101";
	ram(103) <= "0000000000000000000000000000000010000110000000000000000000000000001110000101";
	ram(104) <= "0000000000000000000000000000000011000110000000000000000000000000001110000101";
	ram(105) <= "0000000000000000000000000000000100000110000000000000000000000000001110000101";
	ram(106) <= "0000000000000000000000000000000001000010000000000000000000000000001110000101";
	ram(107) <= "0000000000000000000000000000000010000010000000000000000000000000001110000101";
	ram(108) <= "0000000000000000000000000000000000000000000000000000000000000001000110000100";
	ram(109) <= "0000000000000000000000000000000000000000111000000000000000000000000000000000";
	ram(110) <= "0000000000000000000000000000000001000010000011010000000000000000000000000000";
	ram(111) <= "0000000000000000000000000000000000000000000000000000000000000001001001101110";
	ram(112) <= "0000000000000000000000000000000000000000000101010000000000000000000000000000";
	ram(113) <= "0000000000000000000000000000000000000000110001100000000000000000001110000101";
	ram(114) <= "0000000000000111110000000000000000000000000000000000000000000000000000000000";
	ram(115) <= "0000000000000000000000000000000000000100000000000000000000000000001110000101";
	ram(116) <= "1010000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(117) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(118) <= "0000000000000100000000000000000000000000000000000000000010000000000000000000";
	ram(119) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(120) <= "0000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(121) <= "0000000000000000000000000000000000000100000000000000000000000000001110000101";
	ram(122) <= "1010000000000110000000000000000000000000000000001000000000000000000000000000";
	ram(123) <= "0001010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(124) <= "0000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(125) <= "0001100000000000000000000000000000000000000000000000000010000000000000000000";
	ram(126) <= "0000000000000000000000000000010000000000000000000000000000000000001110000101";
	ram(127) <= "0000000000000000000000000000000110000101000000000000000000000000000000000000";
	ram(128) <= "0000000000000000000000000000000100000101000000000000000000000000001110000101";
	ram(129) <= "0000000000000000000000000000000000000000000001110000000000000000001110000101";
	ram(130) <= "0000000000000000000000000000000000000000000000000100000000000000001110000101";
	ram(131) <= "0000000000000000000000000000000000000000000000000010000000000000001110000101";
	ram(132) <= "0000000000000000000000000000000000000000000000000001000000000000000000000000";
	ram(133) <= "0000000000000000000000000000000000000000000000000000000000000001001110000111";
	ram(134) <= "0000000000000000000000000000000000000000000000000000110101000000001110001101";
	ram(135) <= "0000000000000000000000000000000000000000000000000000000000000001010010001001";
	ram(136) <= "0000000000000000000000000000000000000000000000000000111000100000001110001101";
	ram(137) <= "0000000000000000000000000000000000000000000000000000000000000001010110001011";
	ram(138) <= "0000000000000000000000000000000000000000000000000000111100010000001110001101";
	ram(139) <= "0000000000000000000000000000000000000000000000000000000000000001011000000000";
	ram(140) <= "0000000000000000000000000000000000000000000000000000100000000000000000000000";
	ram(141) <= "0000000000000110010100000000000000000000000000000000000000000000000000000000";
	ram(142) <= "1101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(143) <= "0000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(144) <= "1101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(145) <= "0000000000000110100100000000010000000000000000000000000000000000000000000000";
	ram(146) <= "1101100000000000000000000000000000000000000000000000000000000000000000000000";
	ram(147) <= "0000000000000000000100000000010000000000000000000000000000000000000000000000";
	ram(148) <= "1101010000000000000000000000000000000000000000000000000000000000000000000000";
	ram(149) <= "0000000000000000000000000000010000000000000000000000000000000000000000000000";
	ram(150) <= "1110000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(151) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(152) <= "0000000000000100000000000000000000000000000000000000000010000000000000000000";
	ram(153) <= "0001000000000000000000000000000000000000000000000000000000000000000000000000";
	ram(154) <= "0000000000000010000000000000000000000000000000000000000000000000000000000000";
	ram(155) <= "0000000001000000000000000000000000000000000000000000000000000000001100000000";
	
END description;



--00 00 00 00 00 00 00 00		00 00
