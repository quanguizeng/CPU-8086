LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;
USE ieee.Numeric_Std.ALL;

ENTITY ROM IS
	PORT (
		addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- address
		dat_out  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); -- data to write
		clk : IN STD_LOGIC -- clock
	);
END ENTITY ROM;

ARCHITECTURE description OF ROM IS

   TYPE rom_type IS ARRAY (0 TO 1023) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
   SIGNAL rom : rom_type;

BEGIN	
	dat_out <= rom(to_integer(unsigned(addr)));
	
	rom(0) <= "00000000";
rom(1) <= "00000000";
rom(2) <= "00000000";
rom(3) <= "00000000";
rom(4) <= "00000000";
rom(5) <= "00000000";
rom(6) <= "00000000";
rom(7) <= "00000000";
rom(8) <= "00000000";
rom(9) <= "00000000";
rom(10) <= "00000000";
rom(11) <= "00000000";
rom(12) <= "00000000";
rom(13) <= "00000000";
rom(14) <= "00000000";
rom(15) <= "00000000";
rom(16) <= "00000000";
rom(17) <= "00000000";
rom(18) <= "00000000";
rom(19) <= "00000000";
rom(20) <= "00000000";
rom(21) <= "00000000";
rom(22) <= "00000000";
rom(23) <= "00000000";
rom(24) <= "00000000";
rom(25) <= "00000000";
rom(26) <= "00000000";
rom(27) <= "00000000";
rom(28) <= "00000000";
rom(29) <= "00000000";
rom(30) <= "00000000";
rom(31) <= "00000000";
rom(32) <= "00000000";
rom(33) <= "00000000";
rom(34) <= "00000000";
rom(35) <= "00000000";
rom(36) <= "00000000";
rom(37) <= "00000000";
rom(38) <= "00000000";
rom(39) <= "00000000";
rom(40) <= "00000000";
rom(41) <= "00000000";
rom(42) <= "00000000";
rom(43) <= "00000000";
rom(44) <= "00000000";
rom(45) <= "00000000";
rom(46) <= "00000000";
rom(47) <= "00000000";
rom(48) <= "00000000";
rom(49) <= "00000000";
rom(50) <= "00000000";
rom(51) <= "00000000";
rom(52) <= "00000000";
rom(53) <= "00000000";
rom(54) <= "00000000";
rom(55) <= "00000000";
rom(56) <= "00000000";
rom(57) <= "00000000";
rom(58) <= "00000000";
rom(59) <= "00000000";
rom(60) <= "00000000";
rom(61) <= "00000000";
rom(62) <= "00000000";
rom(63) <= "00000000";
rom(64) <= "00000000";
rom(65) <= "00000000";
rom(66) <= "00000000";
rom(67) <= "00000000";
rom(68) <= "00000000";
rom(69) <= "00000000";
rom(70) <= "00000000";
rom(71) <= "00000000";
rom(72) <= "00000000";
rom(73) <= "00000000";
rom(74) <= "00000000";
rom(75) <= "00000000";
rom(76) <= "00000000";
rom(77) <= "00000000";
rom(78) <= "00000000";
rom(79) <= "00000000";
rom(80) <= "00000000";
rom(81) <= "00000000";
rom(82) <= "00000000";
rom(83) <= "00000000";
rom(84) <= "00000000";
rom(85) <= "00000000";
rom(86) <= "00000000";
rom(87) <= "00000000";
rom(88) <= "00000000";
rom(89) <= "00000000";
rom(90) <= "00000000";
rom(91) <= "00000000";
rom(92) <= "00000000";
rom(93) <= "00000000";
rom(94) <= "00000000";
rom(95) <= "00000000";
rom(96) <= "00000000";
rom(97) <= "00000000";
rom(98) <= "00000000";
rom(99) <= "00000000";
rom(100) <= "00000000";
rom(101) <= "00000000";
rom(102) <= "00000000";
rom(103) <= "00000000";
rom(104) <= "00000000";
rom(105) <= "00000000";
rom(106) <= "00000000";
rom(107) <= "00000000";
rom(108) <= "00000000";
rom(109) <= "00000000";
rom(110) <= "00000000";
rom(111) <= "00000000";
rom(112) <= "00000000";
rom(113) <= "00000000";
rom(114) <= "00000000";
rom(115) <= "00000000";
rom(116) <= "00000000";
rom(117) <= "00000000";
rom(118) <= "00000000";
rom(119) <= "00000000";
rom(120) <= "00000000";
rom(121) <= "00000000";
rom(122) <= "00000000";
rom(123) <= "00000000";
rom(124) <= "00000000";
rom(125) <= "00000000";
rom(126) <= "00000000";
rom(127) <= "00000000";
rom(128) <= "00000000";
rom(129) <= "00000000";
rom(130) <= "00000000";
rom(131) <= "00000000";
rom(132) <= "00000000";
rom(133) <= "00000000";
rom(134) <= "00000000";
rom(135) <= "00000000";
rom(136) <= "00000000";
rom(137) <= "00000000";
rom(138) <= "00000000";
rom(139) <= "00000000";
rom(140) <= "00000000";
rom(141) <= "00000000";
rom(142) <= "00000000";
rom(143) <= "00000000";
rom(144) <= "00000000";
rom(145) <= "00000000";
rom(146) <= "00000000";
rom(147) <= "00000000";
rom(148) <= "00000000";
rom(149) <= "00000000";
rom(150) <= "00000000";
rom(151) <= "00000000";
rom(152) <= "00000000";
rom(153) <= "00000000";
rom(154) <= "00000000";
rom(155) <= "00000000";
rom(156) <= "00000000";
rom(157) <= "00000000";
rom(158) <= "00000000";
rom(159) <= "00000000";
rom(160) <= "00000000";
rom(161) <= "00000000";
rom(162) <= "00000000";
rom(163) <= "00000000";
rom(164) <= "00000000";
rom(165) <= "00000000";
rom(166) <= "00000000";
rom(167) <= "00000000";
rom(168) <= "00000000";
rom(169) <= "00000000";
rom(170) <= "00000000";
rom(171) <= "00000000";
rom(172) <= "00000000";
rom(173) <= "00000000";
rom(174) <= "00000000";
rom(175) <= "00000000";
rom(176) <= "00000000";
rom(177) <= "00000000";
rom(178) <= "00000000";
rom(179) <= "00000000";
rom(180) <= "00000000";
rom(181) <= "00000000";
rom(182) <= "00000000";
rom(183) <= "00000000";
rom(184) <= "00000000";
rom(185) <= "00000000";
rom(186) <= "00000000";
rom(187) <= "00000000";
rom(188) <= "00000000";
rom(189) <= "00000000";
rom(190) <= "00000000";
rom(191) <= "00000000";
rom(192) <= "00000000";
rom(193) <= "00000000";
rom(194) <= "00000000";
rom(195) <= "00000000";
rom(196) <= "00000000";
rom(197) <= "00000000";
rom(198) <= "00000000";
rom(199) <= "00000000";
rom(200) <= "00000000";
rom(201) <= "00000000";
rom(202) <= "00000000";
rom(203) <= "00000000";
rom(204) <= "00000000";
rom(205) <= "00000000";
rom(206) <= "00000000";
rom(207) <= "00000000";
rom(208) <= "00000000";
rom(209) <= "00000000";
rom(210) <= "00000000";
rom(211) <= "00000000";
rom(212) <= "00000000";
rom(213) <= "00000000";
rom(214) <= "00000000";
rom(215) <= "00000000";
rom(216) <= "00000000";
rom(217) <= "00000000";
rom(218) <= "00000000";
rom(219) <= "00000000";
rom(220) <= "00000000";
rom(221) <= "00000000";
rom(222) <= "00000000";
rom(223) <= "00000000";
rom(224) <= "00000000";
rom(225) <= "00000000";
rom(226) <= "00000000";
rom(227) <= "00000000";
rom(228) <= "00000000";
rom(229) <= "00000000";
rom(230) <= "00000000";
rom(231) <= "00000000";
rom(232) <= "00000000";
rom(233) <= "00000000";
rom(234) <= "00000000";
rom(235) <= "00000000";
rom(236) <= "00000000";
rom(237) <= "00000000";
rom(238) <= "00000000";
rom(239) <= "00000000";
rom(240) <= "00000000";
rom(241) <= "00000000";
rom(242) <= "00000000";
rom(243) <= "00000000";
rom(244) <= "00000000";
rom(245) <= "00000000";
rom(246) <= "00000000";
rom(247) <= "00000000";
rom(248) <= "00000000";
rom(249) <= "00000000";
rom(250) <= "00000000";
rom(251) <= "00000000";
rom(252) <= "00000000";
rom(253) <= "00000000";
rom(254) <= "00000000";
rom(255) <= "00000000";
rom(256) <= "00000000";
rom(257) <= "00000000";
rom(258) <= "00000000";
rom(259) <= "00000000";
rom(260) <= "00000000";
rom(261) <= "00000000";
rom(262) <= "00000000";
rom(263) <= "00000000";
rom(264) <= "00000000";
rom(265) <= "00000000";
rom(266) <= "00000000";
rom(267) <= "00000000";
rom(268) <= "00000000";
rom(269) <= "00000000";
rom(270) <= "00000000";
rom(271) <= "00000000";
rom(272) <= "00000000";
rom(273) <= "00000000";
rom(274) <= "00000000";
rom(275) <= "00000000";
rom(276) <= "00000000";
rom(277) <= "00000000";
rom(278) <= "00000000";
rom(279) <= "00000000";
rom(280) <= "00000000";
rom(281) <= "00000000";
rom(282) <= "00000000";
rom(283) <= "00000000";
rom(284) <= "00000000";
rom(285) <= "00000000";
rom(286) <= "00000000";
rom(287) <= "00000000";
rom(288) <= "00000000";
rom(289) <= "00000000";
rom(290) <= "00000000";
rom(291) <= "00000000";
rom(292) <= "00000000";
rom(293) <= "00000000";
rom(294) <= "00000000";
rom(295) <= "00000000";
rom(296) <= "00000000";
rom(297) <= "00000000";
rom(298) <= "00000000";
rom(299) <= "00000000";
rom(300) <= "00000000";
rom(301) <= "00000000";
rom(302) <= "00000000";
rom(303) <= "00000000";
rom(304) <= "00000000";
rom(305) <= "00000000";
rom(306) <= "00000000";
rom(307) <= "00000000";
rom(308) <= "00000000";
rom(309) <= "00000000";
rom(310) <= "00000000";
rom(311) <= "00000000";
rom(312) <= "00000000";
rom(313) <= "00000000";
rom(314) <= "00000000";
rom(315) <= "00000000";
rom(316) <= "00000000";
rom(317) <= "00000000";
rom(318) <= "00000000";
rom(319) <= "00000000";
rom(320) <= "00000000";
rom(321) <= "00000000";
rom(322) <= "00000000";
rom(323) <= "00000000";
rom(324) <= "00000000";
rom(325) <= "00000000";
rom(326) <= "00000000";
rom(327) <= "00000000";
rom(328) <= "00000000";
rom(329) <= "00000000";
rom(330) <= "00000000";
rom(331) <= "00000000";
rom(332) <= "00000000";
rom(333) <= "00000000";
rom(334) <= "00000000";
rom(335) <= "00000000";
rom(336) <= "00000000";
rom(337) <= "00000000";
rom(338) <= "00000000";
rom(339) <= "00000000";
rom(340) <= "00000000";
rom(341) <= "00000000";
rom(342) <= "00000000";
rom(343) <= "00000000";
rom(344) <= "00000000";
rom(345) <= "00000000";
rom(346) <= "00000000";
rom(347) <= "00000000";
rom(348) <= "00000000";
rom(349) <= "00000000";
rom(350) <= "00000000";
rom(351) <= "00000000";
rom(352) <= "00000000";
rom(353) <= "00000000";
rom(354) <= "00000000";
rom(355) <= "00000000";
rom(356) <= "00000000";
rom(357) <= "00000000";
rom(358) <= "00000000";
rom(359) <= "00000000";
rom(360) <= "00000000";
rom(361) <= "00000000";
rom(362) <= "00000000";
rom(363) <= "00000000";
rom(364) <= "00000000";
rom(365) <= "00000000";
rom(366) <= "00000000";
rom(367) <= "00000000";
rom(368) <= "00000000";
rom(369) <= "00000000";
rom(370) <= "00000000";
rom(371) <= "00000000";
rom(372) <= "00000000";
rom(373) <= "00000000";
rom(374) <= "00000000";
rom(375) <= "00000000";
rom(376) <= "00000000";
rom(377) <= "00000000";
rom(378) <= "00000000";
rom(379) <= "00000000";
rom(380) <= "00000000";
rom(381) <= "00000000";
rom(382) <= "00000000";
rom(383) <= "00000000";
rom(384) <= "00000000";
rom(385) <= "00000000";
rom(386) <= "00000000";
rom(387) <= "00000000";
rom(388) <= "00000000";
rom(389) <= "00000000";
rom(390) <= "00000000";
rom(391) <= "00000000";
rom(392) <= "00000000";
rom(393) <= "00000000";
rom(394) <= "00000000";
rom(395) <= "00000000";
rom(396) <= "00000000";
rom(397) <= "00000000";
rom(398) <= "00000000";
rom(399) <= "00000000";
rom(400) <= "00000000";
rom(401) <= "00000000";
rom(402) <= "00000000";
rom(403) <= "00000000";
rom(404) <= "00000000";
rom(405) <= "00000000";
rom(406) <= "00000000";
rom(407) <= "00000000";
rom(408) <= "00000000";
rom(409) <= "00000000";
rom(410) <= "00000000";
rom(411) <= "00000000";
rom(412) <= "00000000";
rom(413) <= "00000000";
rom(414) <= "00000000";
rom(415) <= "00000000";
rom(416) <= "00000000";
rom(417) <= "00000000";
rom(418) <= "00000000";
rom(419) <= "00000000";
rom(420) <= "00000000";
rom(421) <= "00000000";
rom(422) <= "00000000";
rom(423) <= "00000000";
rom(424) <= "00000000";
rom(425) <= "00000000";
rom(426) <= "00000000";
rom(427) <= "00000000";
rom(428) <= "00000000";
rom(429) <= "00000000";
rom(430) <= "00000000";
rom(431) <= "00000000";
rom(432) <= "00000000";
rom(433) <= "00000000";
rom(434) <= "00000000";
rom(435) <= "00000000";
rom(436) <= "00000000";
rom(437) <= "00000000";
rom(438) <= "00000000";
rom(439) <= "00000000";
rom(440) <= "00000000";
rom(441) <= "00000000";
rom(442) <= "00000000";
rom(443) <= "00000000";
rom(444) <= "00000000";
rom(445) <= "00000000";
rom(446) <= "00000000";
rom(447) <= "00000000";
rom(448) <= "00000000";
rom(449) <= "00000000";
rom(450) <= "00000000";
rom(451) <= "00000000";
rom(452) <= "00000000";
rom(453) <= "00000000";
rom(454) <= "00000000";
rom(455) <= "00000000";
rom(456) <= "00000000";
rom(457) <= "00000000";
rom(458) <= "00000000";
rom(459) <= "00000000";
rom(460) <= "00000000";
rom(461) <= "00000000";
rom(462) <= "00000000";
rom(463) <= "00000000";
rom(464) <= "00000000";
rom(465) <= "00000000";
rom(466) <= "00000000";
rom(467) <= "00000000";
rom(468) <= "00000000";
rom(469) <= "00000000";
rom(470) <= "00000000";
rom(471) <= "00000000";
rom(472) <= "00000000";
rom(473) <= "00000000";
rom(474) <= "00000000";
rom(475) <= "00000000";
rom(476) <= "00000000";
rom(477) <= "00000000";
rom(478) <= "00000000";
rom(479) <= "00000000";
rom(480) <= "00000000";
rom(481) <= "00000000";
rom(482) <= "00000000";
rom(483) <= "00000000";
rom(484) <= "00000000";
rom(485) <= "00000000";
rom(486) <= "00000000";
rom(487) <= "00000000";
rom(488) <= "00000000";
rom(489) <= "00000000";
rom(490) <= "00000000";
rom(491) <= "00000000";
rom(492) <= "00000000";
rom(493) <= "00000000";
rom(494) <= "00000000";
rom(495) <= "00000000";
rom(496) <= "00000000";
rom(497) <= "00000000";
rom(498) <= "00000000";
rom(499) <= "00000000";
rom(500) <= "00000000";
rom(501) <= "00000000";
rom(502) <= "00000000";
rom(503) <= "00000000";
rom(504) <= "00000000";
rom(505) <= "00000000";
rom(506) <= "00000000";
rom(507) <= "00000000";
rom(508) <= "00000000";
rom(509) <= "00000000";
rom(510) <= "00000000";
rom(511) <= "00000000";
rom(512) <= "11000000";
rom(513) <= "00010000";
rom(514) <= "00000000";
rom(515) <= "11110100";
rom(516) <= "00000011";
rom(517) <= "00000000";
rom(518) <= "11111000";
rom(519) <= "01011010";
rom(520) <= "10010110";
rom(521) <= "00000000";
rom(522) <= "00000000";
rom(523) <= "00000000";
rom(524) <= "00000000";
rom(525) <= "00000000";
rom(526) <= "00000000";
rom(527) <= "00000000";
rom(528) <= "00000000";
rom(529) <= "00000000";
rom(530) <= "00000000";
rom(531) <= "00000000";
rom(532) <= "00000000";
rom(533) <= "00000000";
rom(534) <= "00000000";
rom(535) <= "00000000";
rom(536) <= "00000000";
rom(537) <= "00000000";
rom(538) <= "00000000";
rom(539) <= "00000000";
rom(540) <= "00000000";
rom(541) <= "00000000";
rom(542) <= "00000000";
rom(543) <= "00000000";
rom(544) <= "00000000";
rom(545) <= "00000000";
rom(546) <= "00000000";
rom(547) <= "00000000";
rom(548) <= "00000000";
rom(549) <= "00000000";
rom(550) <= "00000000";
rom(551) <= "00000000";
rom(552) <= "00000000";
rom(553) <= "00000000";
rom(554) <= "00000000";
rom(555) <= "00000000";
rom(556) <= "00000000";
rom(557) <= "00000000";
rom(558) <= "00000000";
rom(559) <= "00000000";
rom(560) <= "00000000";
rom(561) <= "00000000";
rom(562) <= "00000000";
rom(563) <= "00000000";
rom(564) <= "00000000";
rom(565) <= "00000000";
rom(566) <= "00000000";
rom(567) <= "00000000";
rom(568) <= "00000000";
rom(569) <= "00000000";
rom(570) <= "00000000";
rom(571) <= "00000000";
rom(572) <= "00000000";
rom(573) <= "00000000";
rom(574) <= "00000000";
rom(575) <= "00000000";
rom(576) <= "00000000";
rom(577) <= "00000000";
rom(578) <= "00000000";
rom(579) <= "00000000";
rom(580) <= "00000000";
rom(581) <= "00000000";
rom(582) <= "00000000";
rom(583) <= "00000000";
rom(584) <= "00000000";
rom(585) <= "00000000";
rom(586) <= "00000000";
rom(587) <= "00000000";
rom(588) <= "00000000";
rom(589) <= "00000000";
rom(590) <= "00000000";
rom(591) <= "00000000";
rom(592) <= "00000000";
rom(593) <= "00000000";
rom(594) <= "00000000";
rom(595) <= "00000000";
rom(596) <= "00000000";
rom(597) <= "00000000";
rom(598) <= "00000000";
rom(599) <= "00000000";
rom(600) <= "00000000";
rom(601) <= "00000000";
rom(602) <= "00000000";
rom(603) <= "00000000";
rom(604) <= "00000000";
rom(605) <= "00000000";
rom(606) <= "00000000";
rom(607) <= "00000000";
rom(608) <= "00000000";
rom(609) <= "00000000";
rom(610) <= "00000000";
rom(611) <= "00000000";
rom(612) <= "00000000";
rom(613) <= "00000000";
rom(614) <= "00000000";
rom(615) <= "00000000";
rom(616) <= "00000000";
rom(617) <= "00000000";
rom(618) <= "00000000";
rom(619) <= "00000000";
rom(620) <= "00000000";
rom(621) <= "00000000";
rom(622) <= "00000000";
rom(623) <= "00000000";
rom(624) <= "00000000";
rom(625) <= "00000000";
rom(626) <= "00000000";
rom(627) <= "00000000";
rom(628) <= "00000000";
rom(629) <= "00000000";
rom(630) <= "00000000";
rom(631) <= "00000000";
rom(632) <= "00000000";
rom(633) <= "00000000";
rom(634) <= "00000000";
rom(635) <= "00000000";
rom(636) <= "00000000";
rom(637) <= "00000000";
rom(638) <= "00000000";
rom(639) <= "00000000";
rom(640) <= "00000000";
rom(641) <= "00000000";
rom(642) <= "00000000";
rom(643) <= "00000000";
rom(644) <= "00000000";
rom(645) <= "00000000";
rom(646) <= "00000000";
rom(647) <= "00000000";
rom(648) <= "00000000";
rom(649) <= "00000000";
rom(650) <= "00000000";
rom(651) <= "00000000";
rom(652) <= "00000000";
rom(653) <= "00000000";
rom(654) <= "00000000";
rom(655) <= "00000000";
rom(656) <= "00000000";
rom(657) <= "00000000";
rom(658) <= "00000000";
rom(659) <= "00000000";
rom(660) <= "00000000";
rom(661) <= "00000000";
rom(662) <= "00000000";
rom(663) <= "00000000";
rom(664) <= "00000000";
rom(665) <= "00000000";
rom(666) <= "00000000";
rom(667) <= "00000000";
rom(668) <= "00000000";
rom(669) <= "00000000";
rom(670) <= "00000000";
rom(671) <= "00000000";
rom(672) <= "00000000";
rom(673) <= "00000000";
rom(674) <= "00000000";
rom(675) <= "00000000";
rom(676) <= "00000000";
rom(677) <= "00000000";
rom(678) <= "00000000";
rom(679) <= "00000000";
rom(680) <= "00000000";
rom(681) <= "00000000";
rom(682) <= "00000000";
rom(683) <= "00000000";
rom(684) <= "00000000";
rom(685) <= "00000000";
rom(686) <= "00000000";
rom(687) <= "00000000";
rom(688) <= "00000000";
rom(689) <= "00000000";
rom(690) <= "00000000";
rom(691) <= "00000000";
rom(692) <= "00000000";
rom(693) <= "00000000";
rom(694) <= "00000000";
rom(695) <= "00000000";
rom(696) <= "00000000";
rom(697) <= "00000000";
rom(698) <= "00000000";
rom(699) <= "00000000";
rom(700) <= "00000000";
rom(701) <= "00000000";
rom(702) <= "00000000";
rom(703) <= "00000000";
rom(704) <= "00000000";
rom(705) <= "00000000";
rom(706) <= "00000000";
rom(707) <= "00000000";
rom(708) <= "00000000";
rom(709) <= "00000000";
rom(710) <= "00000000";
rom(711) <= "00000000";
rom(712) <= "00000000";
rom(713) <= "00000000";
rom(714) <= "00000000";
rom(715) <= "00000000";
rom(716) <= "00000000";
rom(717) <= "00000000";
rom(718) <= "00000000";
rom(719) <= "00000000";
rom(720) <= "00000000";
rom(721) <= "00000000";
rom(722) <= "00000000";
rom(723) <= "00000000";
rom(724) <= "00000000";
rom(725) <= "00000000";
rom(726) <= "00000000";
rom(727) <= "00000000";
rom(728) <= "00000000";
rom(729) <= "00000000";
rom(730) <= "00000000";
rom(731) <= "00000000";
rom(732) <= "00000000";
rom(733) <= "00000000";
rom(734) <= "00000000";
rom(735) <= "00000000";
rom(736) <= "00000000";
rom(737) <= "00000000";
rom(738) <= "00000000";
rom(739) <= "00000000";
rom(740) <= "00000000";
rom(741) <= "00000000";
rom(742) <= "00000000";
rom(743) <= "00000000";
rom(744) <= "00000000";
rom(745) <= "00000000";
rom(746) <= "00000000";
rom(747) <= "00000000";
rom(748) <= "00000000";
rom(749) <= "00000000";
rom(750) <= "00000000";
rom(751) <= "00000000";
rom(752) <= "00000000";
rom(753) <= "00000000";
rom(754) <= "00000000";
rom(755) <= "00000000";
rom(756) <= "00000000";
rom(757) <= "00000000";
rom(758) <= "00000000";
rom(759) <= "00000000";
rom(760) <= "00000000";
rom(761) <= "00000000";
rom(762) <= "00000000";
rom(763) <= "00000000";
rom(764) <= "00000000";
rom(765) <= "00000000";
rom(766) <= "00000000";
rom(767) <= "00000000";
rom(768) <= "00000000";
rom(769) <= "00000000";
rom(770) <= "00000000";
rom(771) <= "00000000";
rom(772) <= "00000000";
rom(773) <= "00000000";
rom(774) <= "00000000";
rom(775) <= "00000000";
rom(776) <= "00000000";
rom(777) <= "00000000";
rom(778) <= "00000000";
rom(779) <= "00000000";
rom(780) <= "00000000";
rom(781) <= "00000000";
rom(782) <= "00000000";
rom(783) <= "00000000";
rom(784) <= "00000000";
rom(785) <= "00000000";
rom(786) <= "00000000";
rom(787) <= "00000000";
rom(788) <= "00000000";
rom(789) <= "00000000";
rom(790) <= "00000000";
rom(791) <= "00000000";
rom(792) <= "00000000";
rom(793) <= "00000000";
rom(794) <= "00000000";
rom(795) <= "00000000";
rom(796) <= "00000000";
rom(797) <= "00000000";
rom(798) <= "00000000";
rom(799) <= "00000000";
rom(800) <= "00000000";
rom(801) <= "00000000";
rom(802) <= "00000000";
rom(803) <= "00000000";
rom(804) <= "00000000";
rom(805) <= "00000000";
rom(806) <= "00000000";
rom(807) <= "00000000";
rom(808) <= "00000000";
rom(809) <= "00000000";
rom(810) <= "00000000";
rom(811) <= "00000000";
rom(812) <= "00000000";
rom(813) <= "00000000";
rom(814) <= "00000000";
rom(815) <= "00000000";
rom(816) <= "00000000";
rom(817) <= "00000000";
rom(818) <= "00000000";
rom(819) <= "00000000";
rom(820) <= "00000000";
rom(821) <= "00000000";
rom(822) <= "00000000";
rom(823) <= "00000000";
rom(824) <= "00000000";
rom(825) <= "00000000";
rom(826) <= "00000000";
rom(827) <= "00000000";
rom(828) <= "00000000";
rom(829) <= "00000000";
rom(830) <= "00000000";
rom(831) <= "00000000";
rom(832) <= "00000000";
rom(833) <= "00000000";
rom(834) <= "00000000";
rom(835) <= "00000000";
rom(836) <= "00000000";
rom(837) <= "00000000";
rom(838) <= "00000000";
rom(839) <= "00000000";
rom(840) <= "00000000";
rom(841) <= "00000000";
rom(842) <= "00000000";
rom(843) <= "00000000";
rom(844) <= "00000000";
rom(845) <= "00000000";
rom(846) <= "00000000";
rom(847) <= "00000000";
rom(848) <= "00000000";
rom(849) <= "00000000";
rom(850) <= "00000000";
rom(851) <= "00000000";
rom(852) <= "00000000";
rom(853) <= "00000000";
rom(854) <= "00000000";
rom(855) <= "00000000";
rom(856) <= "00000000";
rom(857) <= "00000000";
rom(858) <= "00000000";
rom(859) <= "00000000";
rom(860) <= "00000000";
rom(861) <= "00000000";
rom(862) <= "00000000";
rom(863) <= "00000000";
rom(864) <= "00000000";
rom(865) <= "00000000";
rom(866) <= "00000000";
rom(867) <= "00000000";
rom(868) <= "00000000";
rom(869) <= "00000000";
rom(870) <= "00000000";
rom(871) <= "00000000";
rom(872) <= "00000000";
rom(873) <= "00000000";
rom(874) <= "00000000";
rom(875) <= "00000000";
rom(876) <= "00000000";
rom(877) <= "00000000";
rom(878) <= "00000000";
rom(879) <= "00000000";
rom(880) <= "00000000";
rom(881) <= "00000000";
rom(882) <= "00000000";
rom(883) <= "00000000";
rom(884) <= "00000000";
rom(885) <= "00000000";
rom(886) <= "00000000";
rom(887) <= "00000000";
rom(888) <= "00000000";
rom(889) <= "00000000";
rom(890) <= "00000000";
rom(891) <= "00000000";
rom(892) <= "00000000";
rom(893) <= "00000000";
rom(894) <= "00000000";
rom(895) <= "00000000";
rom(896) <= "00000000";
rom(897) <= "00000000";
rom(898) <= "00000000";
rom(899) <= "00000000";
rom(900) <= "00000000";
rom(901) <= "00000000";
rom(902) <= "00000000";
rom(903) <= "00000000";
rom(904) <= "00000000";
rom(905) <= "00000000";
rom(906) <= "00000000";
rom(907) <= "00000000";
rom(908) <= "00000000";
rom(909) <= "00000000";
rom(910) <= "00000000";
rom(911) <= "00000000";
rom(912) <= "00000000";
rom(913) <= "00000000";
rom(914) <= "00000000";
rom(915) <= "00000000";
rom(916) <= "00000000";
rom(917) <= "00000000";
rom(918) <= "00000000";
rom(919) <= "00000000";
rom(920) <= "00000000";
rom(921) <= "00000000";
rom(922) <= "00000000";
rom(923) <= "00000000";
rom(924) <= "00000000";
rom(925) <= "00000000";
rom(926) <= "00000000";
rom(927) <= "00000000";
rom(928) <= "00000000";
rom(929) <= "00000000";
rom(930) <= "00000000";
rom(931) <= "00000000";
rom(932) <= "00000000";
rom(933) <= "00000000";
rom(934) <= "00000000";
rom(935) <= "00000000";
rom(936) <= "00000000";
rom(937) <= "00000000";
rom(938) <= "00000000";
rom(939) <= "00000000";
rom(940) <= "00000000";
rom(941) <= "00000000";
rom(942) <= "00000000";
rom(943) <= "00000000";
rom(944) <= "00000000";
rom(945) <= "00000000";
rom(946) <= "00000000";
rom(947) <= "00000000";
rom(948) <= "00000000";
rom(949) <= "00000000";
rom(950) <= "00000000";
rom(951) <= "00000000";
rom(952) <= "00000000";
rom(953) <= "00000000";
rom(954) <= "00000000";
rom(955) <= "00000000";
rom(956) <= "00000000";
rom(957) <= "00000000";
rom(958) <= "00000000";
rom(959) <= "00000000";
rom(960) <= "00000000";
rom(961) <= "00000000";
rom(962) <= "00000000";
rom(963) <= "00000000";
rom(964) <= "00000000";
rom(965) <= "00000000";
rom(966) <= "00000000";
rom(967) <= "00000000";
rom(968) <= "00000000";
rom(969) <= "00000000";
rom(970) <= "00000000";
rom(971) <= "00000000";
rom(972) <= "00000000";
rom(973) <= "00000000";
rom(974) <= "00000000";
rom(975) <= "00000000";
rom(976) <= "00000000";
rom(977) <= "00000000";
rom(978) <= "00000000";
rom(979) <= "00000000";
rom(980) <= "00000000";
rom(981) <= "00000000";
rom(982) <= "00000000";
rom(983) <= "00000000";
rom(984) <= "00000000";
rom(985) <= "00000000";
rom(986) <= "00000000";
rom(987) <= "00000000";
rom(988) <= "00000000";
rom(989) <= "00000000";
rom(990) <= "00000000";
rom(991) <= "00000000";
rom(992) <= "00000000";
rom(993) <= "00000000";
rom(994) <= "00000000";
rom(995) <= "00000000";
rom(996) <= "00000000";
rom(997) <= "00000000";
rom(998) <= "00000000";
rom(999) <= "00000000";
rom(1000) <= "00000000";
rom(1001) <= "00000000";
rom(1002) <= "00000000";
rom(1003) <= "00000000";
rom(1004) <= "00000000";
rom(1005) <= "00000000";
rom(1006) <= "00000000";
rom(1007) <= "00000000";
rom(1008) <= "00000000";
rom(1009) <= "00000000";
rom(1010) <= "00000000";
rom(1011) <= "00000000";
rom(1012) <= "00000000";
rom(1013) <= "00000000";
rom(1014) <= "00000000";
rom(1015) <= "00000000";
rom(1016) <= "00000000";
rom(1017) <= "00000000";
rom(1018) <= "00000000";
rom(1019) <= "00000000";
rom(1020) <= "00000000";
rom(1021) <= "00000000";
rom(1022) <= "00000000";
rom(1023) <= "00000000";

	
END description;
